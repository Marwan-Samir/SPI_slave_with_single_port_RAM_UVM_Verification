interface wrapper_ref_if(clk);

  input clk;
  logic rst_n;
  logic MOSI_ref;
  logic MISO_ref;
  logic SS_n_ref;

endinterface
