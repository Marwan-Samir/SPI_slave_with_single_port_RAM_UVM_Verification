interface wrapper_if(clk);

  input clk;
  logic rst_n;
  logic MOSI;
  logic MISO;
  logic SS_n;

endinterface 
